/*
class slave_seqs extends uvm_sequence#(slave_xtn);

   `uvm_component_utils(slave_seqs)
    extern function new(string name ="slave_seqs", uvm_component parent);
endclass


//-------------------------Constructor-----------------------------//
	function slave_seqs::new(string name = "slave_seqs",uvm_component parent);
	   super.new(name,parent);
  endfunction
*/